import test::* ;
import test2::* ;


module test3 #()();


initial begin
    test_task();
end

endmodule