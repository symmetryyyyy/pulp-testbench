package test;

task test_task;

  $display("1");

endtask

endpackage