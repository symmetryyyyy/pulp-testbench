package test2;

task test_task;

  $display("2");

endtask

endpackage